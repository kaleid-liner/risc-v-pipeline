
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h2d2aa557;
    ram_cell[       1] = 32'h0;  // 32'hb341e718;
    ram_cell[       2] = 32'h0;  // 32'hc2967490;
    ram_cell[       3] = 32'h0;  // 32'h6e0b3df7;
    ram_cell[       4] = 32'h0;  // 32'h4dd4859d;
    ram_cell[       5] = 32'h0;  // 32'hbb5bf19e;
    ram_cell[       6] = 32'h0;  // 32'h46cba0a1;
    ram_cell[       7] = 32'h0;  // 32'h45def5fa;
    ram_cell[       8] = 32'h0;  // 32'h7adcb337;
    ram_cell[       9] = 32'h0;  // 32'h94391aca;
    ram_cell[      10] = 32'h0;  // 32'h5aea464e;
    ram_cell[      11] = 32'h0;  // 32'h66be76a8;
    ram_cell[      12] = 32'h0;  // 32'h7910a038;
    ram_cell[      13] = 32'h0;  // 32'h4f44d449;
    ram_cell[      14] = 32'h0;  // 32'hee061fb7;
    ram_cell[      15] = 32'h0;  // 32'h898476cb;
    ram_cell[      16] = 32'h0;  // 32'haa53e92c;
    ram_cell[      17] = 32'h0;  // 32'h6d9fdc32;
    ram_cell[      18] = 32'h0;  // 32'h6ea48d02;
    ram_cell[      19] = 32'h0;  // 32'h6746da76;
    ram_cell[      20] = 32'h0;  // 32'hb2b8fa1c;
    ram_cell[      21] = 32'h0;  // 32'hca47cffe;
    ram_cell[      22] = 32'h0;  // 32'hb5f4a153;
    ram_cell[      23] = 32'h0;  // 32'h9ea3b2c8;
    ram_cell[      24] = 32'h0;  // 32'h2f1135a8;
    ram_cell[      25] = 32'h0;  // 32'h9a1f9d45;
    ram_cell[      26] = 32'h0;  // 32'h9b80e54d;
    ram_cell[      27] = 32'h0;  // 32'h75157719;
    ram_cell[      28] = 32'h0;  // 32'hbbe7ba34;
    ram_cell[      29] = 32'h0;  // 32'h5033a7c6;
    ram_cell[      30] = 32'h0;  // 32'h7d2db0ff;
    ram_cell[      31] = 32'h0;  // 32'he8d5b5f2;
    ram_cell[      32] = 32'h0;  // 32'h41299f1c;
    ram_cell[      33] = 32'h0;  // 32'h12766052;
    ram_cell[      34] = 32'h0;  // 32'h3028ae40;
    ram_cell[      35] = 32'h0;  // 32'h19fdd639;
    ram_cell[      36] = 32'h0;  // 32'h9ac2e5bb;
    ram_cell[      37] = 32'h0;  // 32'h16fefefd;
    ram_cell[      38] = 32'h0;  // 32'h35c4c5c0;
    ram_cell[      39] = 32'h0;  // 32'h4418d78b;
    ram_cell[      40] = 32'h0;  // 32'h73378244;
    ram_cell[      41] = 32'h0;  // 32'hf2473b0c;
    ram_cell[      42] = 32'h0;  // 32'hc5281154;
    ram_cell[      43] = 32'h0;  // 32'he2850af5;
    ram_cell[      44] = 32'h0;  // 32'h02222bf1;
    ram_cell[      45] = 32'h0;  // 32'h168c78fd;
    ram_cell[      46] = 32'h0;  // 32'h12c5e6ef;
    ram_cell[      47] = 32'h0;  // 32'h80516c0d;
    ram_cell[      48] = 32'h0;  // 32'ha62a7bb6;
    ram_cell[      49] = 32'h0;  // 32'h23505aea;
    ram_cell[      50] = 32'h0;  // 32'hf9648161;
    ram_cell[      51] = 32'h0;  // 32'h864b0ce6;
    ram_cell[      52] = 32'h0;  // 32'h414db7d2;
    ram_cell[      53] = 32'h0;  // 32'h7c4d63e6;
    ram_cell[      54] = 32'h0;  // 32'h381183d6;
    ram_cell[      55] = 32'h0;  // 32'h95050ca3;
    ram_cell[      56] = 32'h0;  // 32'hde6fb327;
    ram_cell[      57] = 32'h0;  // 32'hcfca9fdb;
    ram_cell[      58] = 32'h0;  // 32'he4064a17;
    ram_cell[      59] = 32'h0;  // 32'hdc0b1cec;
    ram_cell[      60] = 32'h0;  // 32'h4d7b5832;
    ram_cell[      61] = 32'h0;  // 32'h83563878;
    ram_cell[      62] = 32'h0;  // 32'h8c6845eb;
    ram_cell[      63] = 32'h0;  // 32'h4f42af59;
    ram_cell[      64] = 32'h0;  // 32'hcb78510d;
    ram_cell[      65] = 32'h0;  // 32'h1fbb84a4;
    ram_cell[      66] = 32'h0;  // 32'h14203741;
    ram_cell[      67] = 32'h0;  // 32'h1bc8b1a2;
    ram_cell[      68] = 32'h0;  // 32'hcea90c9a;
    ram_cell[      69] = 32'h0;  // 32'h29663ef5;
    ram_cell[      70] = 32'h0;  // 32'h7245afcc;
    ram_cell[      71] = 32'h0;  // 32'h93b4a7bb;
    ram_cell[      72] = 32'h0;  // 32'h146913b7;
    ram_cell[      73] = 32'h0;  // 32'h6d3aa7e4;
    ram_cell[      74] = 32'h0;  // 32'h144ef6d7;
    ram_cell[      75] = 32'h0;  // 32'h71b677db;
    ram_cell[      76] = 32'h0;  // 32'h3c0f4667;
    ram_cell[      77] = 32'h0;  // 32'h94010cde;
    ram_cell[      78] = 32'h0;  // 32'h60b430ee;
    ram_cell[      79] = 32'h0;  // 32'h004a4a1a;
    ram_cell[      80] = 32'h0;  // 32'hb5fce0a3;
    ram_cell[      81] = 32'h0;  // 32'hd3219e2c;
    ram_cell[      82] = 32'h0;  // 32'hee8e831e;
    ram_cell[      83] = 32'h0;  // 32'haba0449b;
    ram_cell[      84] = 32'h0;  // 32'h2106264a;
    ram_cell[      85] = 32'h0;  // 32'h111f78ff;
    ram_cell[      86] = 32'h0;  // 32'h85ab45b1;
    ram_cell[      87] = 32'h0;  // 32'h1baa6754;
    ram_cell[      88] = 32'h0;  // 32'h814b915c;
    ram_cell[      89] = 32'h0;  // 32'h02264444;
    ram_cell[      90] = 32'h0;  // 32'h43917e98;
    ram_cell[      91] = 32'h0;  // 32'he8c49432;
    ram_cell[      92] = 32'h0;  // 32'he4b8553d;
    ram_cell[      93] = 32'h0;  // 32'hcef85e6d;
    ram_cell[      94] = 32'h0;  // 32'hc37e3a3a;
    ram_cell[      95] = 32'h0;  // 32'h54fab544;
    ram_cell[      96] = 32'h0;  // 32'ha83583d2;
    ram_cell[      97] = 32'h0;  // 32'h1021af69;
    ram_cell[      98] = 32'h0;  // 32'he53a89db;
    ram_cell[      99] = 32'h0;  // 32'h45bcf912;
    ram_cell[     100] = 32'h0;  // 32'hd29ea62b;
    ram_cell[     101] = 32'h0;  // 32'hac843bdd;
    ram_cell[     102] = 32'h0;  // 32'hff299143;
    ram_cell[     103] = 32'h0;  // 32'h0afe6c30;
    ram_cell[     104] = 32'h0;  // 32'h506893c9;
    ram_cell[     105] = 32'h0;  // 32'h5661ac31;
    ram_cell[     106] = 32'h0;  // 32'he6cea487;
    ram_cell[     107] = 32'h0;  // 32'h49b65f8c;
    ram_cell[     108] = 32'h0;  // 32'h4f865e6d;
    ram_cell[     109] = 32'h0;  // 32'h1674cbef;
    ram_cell[     110] = 32'h0;  // 32'h122d95ab;
    ram_cell[     111] = 32'h0;  // 32'h8d1a7084;
    ram_cell[     112] = 32'h0;  // 32'hb28d87d5;
    ram_cell[     113] = 32'h0;  // 32'hbdf80115;
    ram_cell[     114] = 32'h0;  // 32'h1f51fd32;
    ram_cell[     115] = 32'h0;  // 32'h9ec57e59;
    ram_cell[     116] = 32'h0;  // 32'h250fd55b;
    ram_cell[     117] = 32'h0;  // 32'he5b13310;
    ram_cell[     118] = 32'h0;  // 32'h61245f2a;
    ram_cell[     119] = 32'h0;  // 32'h35bafa02;
    ram_cell[     120] = 32'h0;  // 32'h219e675e;
    ram_cell[     121] = 32'h0;  // 32'hef75086e;
    ram_cell[     122] = 32'h0;  // 32'hdb5dc9de;
    ram_cell[     123] = 32'h0;  // 32'h17b6243f;
    ram_cell[     124] = 32'h0;  // 32'h8638126b;
    ram_cell[     125] = 32'h0;  // 32'h11a689b7;
    ram_cell[     126] = 32'h0;  // 32'h31a8615c;
    ram_cell[     127] = 32'h0;  // 32'hf8fbe8c2;
    ram_cell[     128] = 32'h0;  // 32'hc39d9d73;
    ram_cell[     129] = 32'h0;  // 32'hfe1b35b4;
    ram_cell[     130] = 32'h0;  // 32'h7bd5e8a4;
    ram_cell[     131] = 32'h0;  // 32'h88c9cfd1;
    ram_cell[     132] = 32'h0;  // 32'hb7408940;
    ram_cell[     133] = 32'h0;  // 32'h6d20f507;
    ram_cell[     134] = 32'h0;  // 32'h3f0fe18c;
    ram_cell[     135] = 32'h0;  // 32'hd32636d5;
    ram_cell[     136] = 32'h0;  // 32'h0755dc99;
    ram_cell[     137] = 32'h0;  // 32'h7a0c20db;
    ram_cell[     138] = 32'h0;  // 32'hcd9c7355;
    ram_cell[     139] = 32'h0;  // 32'h95e2b04f;
    ram_cell[     140] = 32'h0;  // 32'h8abc10a5;
    ram_cell[     141] = 32'h0;  // 32'h94569c24;
    ram_cell[     142] = 32'h0;  // 32'hb96211dc;
    ram_cell[     143] = 32'h0;  // 32'h9eecb31b;
    ram_cell[     144] = 32'h0;  // 32'hf84666f1;
    ram_cell[     145] = 32'h0;  // 32'h76b41adf;
    ram_cell[     146] = 32'h0;  // 32'h464fdfe9;
    ram_cell[     147] = 32'h0;  // 32'h5fa2289d;
    ram_cell[     148] = 32'h0;  // 32'hd41c74a6;
    ram_cell[     149] = 32'h0;  // 32'h0bae7e76;
    ram_cell[     150] = 32'h0;  // 32'he6b14558;
    ram_cell[     151] = 32'h0;  // 32'h18f0f1f7;
    ram_cell[     152] = 32'h0;  // 32'h8148d770;
    ram_cell[     153] = 32'h0;  // 32'h4c204552;
    ram_cell[     154] = 32'h0;  // 32'hef1eaedf;
    ram_cell[     155] = 32'h0;  // 32'h03e32796;
    ram_cell[     156] = 32'h0;  // 32'hb9d310b8;
    ram_cell[     157] = 32'h0;  // 32'h2eb0cd73;
    ram_cell[     158] = 32'h0;  // 32'hb89d970c;
    ram_cell[     159] = 32'h0;  // 32'hd78dd1b7;
    ram_cell[     160] = 32'h0;  // 32'hbc46846a;
    ram_cell[     161] = 32'h0;  // 32'hb7340003;
    ram_cell[     162] = 32'h0;  // 32'h49458d57;
    ram_cell[     163] = 32'h0;  // 32'h4a8906f3;
    ram_cell[     164] = 32'h0;  // 32'h43ae422b;
    ram_cell[     165] = 32'h0;  // 32'hff3da4ab;
    ram_cell[     166] = 32'h0;  // 32'h0aa9bc9f;
    ram_cell[     167] = 32'h0;  // 32'h475b96ab;
    ram_cell[     168] = 32'h0;  // 32'h74efd66d;
    ram_cell[     169] = 32'h0;  // 32'hcc948595;
    ram_cell[     170] = 32'h0;  // 32'ha353573f;
    ram_cell[     171] = 32'h0;  // 32'h295161a5;
    ram_cell[     172] = 32'h0;  // 32'h1f8382be;
    ram_cell[     173] = 32'h0;  // 32'hdc3db6ce;
    ram_cell[     174] = 32'h0;  // 32'hd1a44fb5;
    ram_cell[     175] = 32'h0;  // 32'h10750253;
    ram_cell[     176] = 32'h0;  // 32'h8c6c9ca8;
    ram_cell[     177] = 32'h0;  // 32'h526ff4cc;
    ram_cell[     178] = 32'h0;  // 32'h970c9bf5;
    ram_cell[     179] = 32'h0;  // 32'h4f905e89;
    ram_cell[     180] = 32'h0;  // 32'h7f5a3eba;
    ram_cell[     181] = 32'h0;  // 32'hf6b13a8e;
    ram_cell[     182] = 32'h0;  // 32'h74082ea4;
    ram_cell[     183] = 32'h0;  // 32'h860cbe12;
    ram_cell[     184] = 32'h0;  // 32'h80769c0a;
    ram_cell[     185] = 32'h0;  // 32'hdd34ca86;
    ram_cell[     186] = 32'h0;  // 32'h13372431;
    ram_cell[     187] = 32'h0;  // 32'he053a807;
    ram_cell[     188] = 32'h0;  // 32'hc4510236;
    ram_cell[     189] = 32'h0;  // 32'h9626c09d;
    ram_cell[     190] = 32'h0;  // 32'h3bdf4c75;
    ram_cell[     191] = 32'h0;  // 32'h3fc12dd8;
    ram_cell[     192] = 32'h0;  // 32'h6790f876;
    ram_cell[     193] = 32'h0;  // 32'h21073532;
    ram_cell[     194] = 32'h0;  // 32'h2effc724;
    ram_cell[     195] = 32'h0;  // 32'hc77d1e57;
    ram_cell[     196] = 32'h0;  // 32'h96b74c54;
    ram_cell[     197] = 32'h0;  // 32'h7460edaf;
    ram_cell[     198] = 32'h0;  // 32'h34d90672;
    ram_cell[     199] = 32'h0;  // 32'hbdd4428a;
    ram_cell[     200] = 32'h0;  // 32'h96bc2eb7;
    ram_cell[     201] = 32'h0;  // 32'hc3c76d53;
    ram_cell[     202] = 32'h0;  // 32'h16f26e1d;
    ram_cell[     203] = 32'h0;  // 32'h6bdce269;
    ram_cell[     204] = 32'h0;  // 32'h66b705c2;
    ram_cell[     205] = 32'h0;  // 32'ha841f7ef;
    ram_cell[     206] = 32'h0;  // 32'hcb352e35;
    ram_cell[     207] = 32'h0;  // 32'h76681f06;
    ram_cell[     208] = 32'h0;  // 32'h0eeb3eab;
    ram_cell[     209] = 32'h0;  // 32'h9df995b9;
    ram_cell[     210] = 32'h0;  // 32'h1b50d5c2;
    ram_cell[     211] = 32'h0;  // 32'hccf27531;
    ram_cell[     212] = 32'h0;  // 32'h6515e20a;
    ram_cell[     213] = 32'h0;  // 32'h2bcd4591;
    ram_cell[     214] = 32'h0;  // 32'hb3d568a2;
    ram_cell[     215] = 32'h0;  // 32'h877846fa;
    ram_cell[     216] = 32'h0;  // 32'h105bf6a0;
    ram_cell[     217] = 32'h0;  // 32'hd1cdbca7;
    ram_cell[     218] = 32'h0;  // 32'h05be1e1f;
    ram_cell[     219] = 32'h0;  // 32'h0b237b81;
    ram_cell[     220] = 32'h0;  // 32'heef1e125;
    ram_cell[     221] = 32'h0;  // 32'h63cb924a;
    ram_cell[     222] = 32'h0;  // 32'h4ecf4468;
    ram_cell[     223] = 32'h0;  // 32'h3a118c8d;
    ram_cell[     224] = 32'h0;  // 32'h394e3544;
    ram_cell[     225] = 32'h0;  // 32'h698ab76d;
    ram_cell[     226] = 32'h0;  // 32'h1d134d39;
    ram_cell[     227] = 32'h0;  // 32'h4a655578;
    ram_cell[     228] = 32'h0;  // 32'hba594726;
    ram_cell[     229] = 32'h0;  // 32'h8125bd64;
    ram_cell[     230] = 32'h0;  // 32'hd5e4c92f;
    ram_cell[     231] = 32'h0;  // 32'hf83e146c;
    ram_cell[     232] = 32'h0;  // 32'h6c514d0d;
    ram_cell[     233] = 32'h0;  // 32'h2bc10425;
    ram_cell[     234] = 32'h0;  // 32'h4e17e39d;
    ram_cell[     235] = 32'h0;  // 32'hc15b0e03;
    ram_cell[     236] = 32'h0;  // 32'h42efff6c;
    ram_cell[     237] = 32'h0;  // 32'hf85bea96;
    ram_cell[     238] = 32'h0;  // 32'h1b80a2a5;
    ram_cell[     239] = 32'h0;  // 32'h3bc4045c;
    ram_cell[     240] = 32'h0;  // 32'h2c2c04ad;
    ram_cell[     241] = 32'h0;  // 32'h41aec67c;
    ram_cell[     242] = 32'h0;  // 32'ha618b60d;
    ram_cell[     243] = 32'h0;  // 32'h82e0b6c7;
    ram_cell[     244] = 32'h0;  // 32'h23ae997e;
    ram_cell[     245] = 32'h0;  // 32'h2e1a34a3;
    ram_cell[     246] = 32'h0;  // 32'hb977e83c;
    ram_cell[     247] = 32'h0;  // 32'h2228b864;
    ram_cell[     248] = 32'h0;  // 32'he2e16425;
    ram_cell[     249] = 32'h0;  // 32'h65ee3059;
    ram_cell[     250] = 32'h0;  // 32'hfe18a64b;
    ram_cell[     251] = 32'h0;  // 32'h045d322a;
    ram_cell[     252] = 32'h0;  // 32'h6a7018a1;
    ram_cell[     253] = 32'h0;  // 32'h9b24330d;
    ram_cell[     254] = 32'h0;  // 32'hc418548d;
    ram_cell[     255] = 32'h0;  // 32'h8fbb1389;
    // src matrix A
    ram_cell[     256] = 32'hc18f7a83;
    ram_cell[     257] = 32'h40b3d174;
    ram_cell[     258] = 32'h3c70e05b;
    ram_cell[     259] = 32'h33c38ab0;
    ram_cell[     260] = 32'h15ee90b1;
    ram_cell[     261] = 32'hae414990;
    ram_cell[     262] = 32'hf31d5ca8;
    ram_cell[     263] = 32'h7e32cb0a;
    ram_cell[     264] = 32'h492de7fc;
    ram_cell[     265] = 32'h96db6533;
    ram_cell[     266] = 32'h1f3d6613;
    ram_cell[     267] = 32'h31fca566;
    ram_cell[     268] = 32'h80dc3373;
    ram_cell[     269] = 32'h88ed3391;
    ram_cell[     270] = 32'hcc7a20d2;
    ram_cell[     271] = 32'h8611b076;
    ram_cell[     272] = 32'h383a1f28;
    ram_cell[     273] = 32'ha2bb23c0;
    ram_cell[     274] = 32'h9cd73b5e;
    ram_cell[     275] = 32'h37313a20;
    ram_cell[     276] = 32'he156d9e9;
    ram_cell[     277] = 32'h25815deb;
    ram_cell[     278] = 32'h9e765f7c;
    ram_cell[     279] = 32'h79baef84;
    ram_cell[     280] = 32'h0dd94371;
    ram_cell[     281] = 32'had2a18bd;
    ram_cell[     282] = 32'h6f7574e4;
    ram_cell[     283] = 32'hd573671c;
    ram_cell[     284] = 32'h3af339c9;
    ram_cell[     285] = 32'hfc928fcf;
    ram_cell[     286] = 32'h83ad5d63;
    ram_cell[     287] = 32'h1deb4a30;
    ram_cell[     288] = 32'h9b5313bc;
    ram_cell[     289] = 32'h4611103c;
    ram_cell[     290] = 32'h04df6274;
    ram_cell[     291] = 32'h20d3f138;
    ram_cell[     292] = 32'hf5a97dee;
    ram_cell[     293] = 32'hbe723400;
    ram_cell[     294] = 32'hb31dbfae;
    ram_cell[     295] = 32'h81258152;
    ram_cell[     296] = 32'h01dd4021;
    ram_cell[     297] = 32'he84cff11;
    ram_cell[     298] = 32'h05691277;
    ram_cell[     299] = 32'h9f140af6;
    ram_cell[     300] = 32'h63e86455;
    ram_cell[     301] = 32'h01d3d436;
    ram_cell[     302] = 32'h9153ce65;
    ram_cell[     303] = 32'h8d25bc33;
    ram_cell[     304] = 32'hb66da326;
    ram_cell[     305] = 32'hf0bd40dd;
    ram_cell[     306] = 32'hbdb6ab5d;
    ram_cell[     307] = 32'hf4ca1484;
    ram_cell[     308] = 32'h43a8ee3c;
    ram_cell[     309] = 32'hf4794662;
    ram_cell[     310] = 32'hb4dd2f82;
    ram_cell[     311] = 32'h382e13a1;
    ram_cell[     312] = 32'h8cb452d6;
    ram_cell[     313] = 32'h99d90b94;
    ram_cell[     314] = 32'h1ce498dd;
    ram_cell[     315] = 32'ha3e18a14;
    ram_cell[     316] = 32'h9a617567;
    ram_cell[     317] = 32'h797c3889;
    ram_cell[     318] = 32'hd35348a3;
    ram_cell[     319] = 32'haa6cf785;
    ram_cell[     320] = 32'hc8b06718;
    ram_cell[     321] = 32'hb64ba4e9;
    ram_cell[     322] = 32'h59e7a8f1;
    ram_cell[     323] = 32'h75fe0aa9;
    ram_cell[     324] = 32'h74557084;
    ram_cell[     325] = 32'h190c8db6;
    ram_cell[     326] = 32'h23b4a8f5;
    ram_cell[     327] = 32'h404bfda9;
    ram_cell[     328] = 32'hded88782;
    ram_cell[     329] = 32'hafbaf915;
    ram_cell[     330] = 32'hdf674ee8;
    ram_cell[     331] = 32'h5d26850f;
    ram_cell[     332] = 32'h99df86a1;
    ram_cell[     333] = 32'h2b13466f;
    ram_cell[     334] = 32'h2e8943e1;
    ram_cell[     335] = 32'h8d22734c;
    ram_cell[     336] = 32'h6e55c457;
    ram_cell[     337] = 32'hbcf4e8b0;
    ram_cell[     338] = 32'hf35d4850;
    ram_cell[     339] = 32'h977a8db7;
    ram_cell[     340] = 32'h92e471e9;
    ram_cell[     341] = 32'he0f6303b;
    ram_cell[     342] = 32'h96c37078;
    ram_cell[     343] = 32'h4c9bf8df;
    ram_cell[     344] = 32'hef08274d;
    ram_cell[     345] = 32'hb4c8497f;
    ram_cell[     346] = 32'h272d8bac;
    ram_cell[     347] = 32'h7b407fc7;
    ram_cell[     348] = 32'h8a31f1fc;
    ram_cell[     349] = 32'h0fd4ba33;
    ram_cell[     350] = 32'hee5a3ac4;
    ram_cell[     351] = 32'hf3d223fb;
    ram_cell[     352] = 32'hdfa37cdc;
    ram_cell[     353] = 32'h10024871;
    ram_cell[     354] = 32'h138b5fdb;
    ram_cell[     355] = 32'h423b5c7d;
    ram_cell[     356] = 32'hbabbc0e2;
    ram_cell[     357] = 32'hade376b3;
    ram_cell[     358] = 32'h6c8cda76;
    ram_cell[     359] = 32'h11f7a615;
    ram_cell[     360] = 32'h35779dc9;
    ram_cell[     361] = 32'had557e67;
    ram_cell[     362] = 32'hc322245f;
    ram_cell[     363] = 32'h788d8067;
    ram_cell[     364] = 32'hbfd27d3a;
    ram_cell[     365] = 32'h2b031a84;
    ram_cell[     366] = 32'hc3d0f117;
    ram_cell[     367] = 32'h4f171c2c;
    ram_cell[     368] = 32'hc2069127;
    ram_cell[     369] = 32'h29d9b092;
    ram_cell[     370] = 32'h835aeb07;
    ram_cell[     371] = 32'h629c654b;
    ram_cell[     372] = 32'hc65241a8;
    ram_cell[     373] = 32'ha65a2a86;
    ram_cell[     374] = 32'h4eabb838;
    ram_cell[     375] = 32'h5fc30a80;
    ram_cell[     376] = 32'h8debbad1;
    ram_cell[     377] = 32'h7499ad46;
    ram_cell[     378] = 32'h53c22170;
    ram_cell[     379] = 32'h8dfab65e;
    ram_cell[     380] = 32'h19abac31;
    ram_cell[     381] = 32'h018acebc;
    ram_cell[     382] = 32'h42153f15;
    ram_cell[     383] = 32'h38ca174f;
    ram_cell[     384] = 32'h572c26b6;
    ram_cell[     385] = 32'hd53162b1;
    ram_cell[     386] = 32'hc003a517;
    ram_cell[     387] = 32'h03a67dc5;
    ram_cell[     388] = 32'h82aa7d20;
    ram_cell[     389] = 32'h1d5712e4;
    ram_cell[     390] = 32'hf29d97ee;
    ram_cell[     391] = 32'h71e99479;
    ram_cell[     392] = 32'hb76a9032;
    ram_cell[     393] = 32'h63e5fa0a;
    ram_cell[     394] = 32'h09a97e3e;
    ram_cell[     395] = 32'hf5c09ad5;
    ram_cell[     396] = 32'h4480bf45;
    ram_cell[     397] = 32'h240e27ae;
    ram_cell[     398] = 32'hdecc96a4;
    ram_cell[     399] = 32'hf848c008;
    ram_cell[     400] = 32'h146fc10e;
    ram_cell[     401] = 32'h953bcf37;
    ram_cell[     402] = 32'he14d9123;
    ram_cell[     403] = 32'h533bc932;
    ram_cell[     404] = 32'h3a2f9439;
    ram_cell[     405] = 32'h8a542071;
    ram_cell[     406] = 32'h0340ef0f;
    ram_cell[     407] = 32'h569ba953;
    ram_cell[     408] = 32'hcfae608d;
    ram_cell[     409] = 32'h37c85a1a;
    ram_cell[     410] = 32'h80684eaa;
    ram_cell[     411] = 32'hcd55e788;
    ram_cell[     412] = 32'hd61b36a7;
    ram_cell[     413] = 32'hb7b76eb6;
    ram_cell[     414] = 32'had64fc17;
    ram_cell[     415] = 32'hdbf930b2;
    ram_cell[     416] = 32'h45271124;
    ram_cell[     417] = 32'h87aec072;
    ram_cell[     418] = 32'h384c7fe1;
    ram_cell[     419] = 32'haf3c49cf;
    ram_cell[     420] = 32'ha6a506d1;
    ram_cell[     421] = 32'h23444520;
    ram_cell[     422] = 32'hd15a63a9;
    ram_cell[     423] = 32'h4fd59e49;
    ram_cell[     424] = 32'h7d6e8d09;
    ram_cell[     425] = 32'h65a3a74c;
    ram_cell[     426] = 32'hb0d64ccc;
    ram_cell[     427] = 32'hbe171b5d;
    ram_cell[     428] = 32'hbafce398;
    ram_cell[     429] = 32'h3109a4e2;
    ram_cell[     430] = 32'h1b987dd8;
    ram_cell[     431] = 32'hcdbbd7df;
    ram_cell[     432] = 32'hf0feab7e;
    ram_cell[     433] = 32'h928f5557;
    ram_cell[     434] = 32'h7b43e7a3;
    ram_cell[     435] = 32'h1ce90383;
    ram_cell[     436] = 32'h49b30370;
    ram_cell[     437] = 32'he1316f01;
    ram_cell[     438] = 32'h30f8c410;
    ram_cell[     439] = 32'h2cfaef98;
    ram_cell[     440] = 32'ha97ba42f;
    ram_cell[     441] = 32'h6df17baf;
    ram_cell[     442] = 32'h88a94f99;
    ram_cell[     443] = 32'h6ce66c78;
    ram_cell[     444] = 32'h66615584;
    ram_cell[     445] = 32'h6428859d;
    ram_cell[     446] = 32'h2f92f2e2;
    ram_cell[     447] = 32'h09645f73;
    ram_cell[     448] = 32'hb8369b4b;
    ram_cell[     449] = 32'h7a7bdafb;
    ram_cell[     450] = 32'h5ef4c1e7;
    ram_cell[     451] = 32'hc06ce783;
    ram_cell[     452] = 32'h82b9caef;
    ram_cell[     453] = 32'hc31845e8;
    ram_cell[     454] = 32'hfd7a71dc;
    ram_cell[     455] = 32'h21221988;
    ram_cell[     456] = 32'h09d17c5a;
    ram_cell[     457] = 32'h0f6ac7da;
    ram_cell[     458] = 32'hf146b0b8;
    ram_cell[     459] = 32'h1057c958;
    ram_cell[     460] = 32'ha3f289a6;
    ram_cell[     461] = 32'h4cfbc01e;
    ram_cell[     462] = 32'h1f710c2e;
    ram_cell[     463] = 32'he6657a72;
    ram_cell[     464] = 32'h9781731c;
    ram_cell[     465] = 32'h536823b9;
    ram_cell[     466] = 32'h332e1ec7;
    ram_cell[     467] = 32'h0f1fb58b;
    ram_cell[     468] = 32'h2c2c7026;
    ram_cell[     469] = 32'hb8cee2ac;
    ram_cell[     470] = 32'he46524e3;
    ram_cell[     471] = 32'h64b0f622;
    ram_cell[     472] = 32'h2e75d4ea;
    ram_cell[     473] = 32'he7453476;
    ram_cell[     474] = 32'h31249a04;
    ram_cell[     475] = 32'h8c893a70;
    ram_cell[     476] = 32'h2233e052;
    ram_cell[     477] = 32'h4041ab1e;
    ram_cell[     478] = 32'h93c4d01e;
    ram_cell[     479] = 32'h0a66481f;
    ram_cell[     480] = 32'he32fa0b1;
    ram_cell[     481] = 32'h19aa83b5;
    ram_cell[     482] = 32'h3c28a5da;
    ram_cell[     483] = 32'h4f401035;
    ram_cell[     484] = 32'h87d08764;
    ram_cell[     485] = 32'h3f1acaf0;
    ram_cell[     486] = 32'h8b56d432;
    ram_cell[     487] = 32'he148e972;
    ram_cell[     488] = 32'h8ef96ef1;
    ram_cell[     489] = 32'hee18b2da;
    ram_cell[     490] = 32'h4a486566;
    ram_cell[     491] = 32'h6867e2ca;
    ram_cell[     492] = 32'ha7350651;
    ram_cell[     493] = 32'h3e5d7fc8;
    ram_cell[     494] = 32'he455012a;
    ram_cell[     495] = 32'h6c179621;
    ram_cell[     496] = 32'h9020bf39;
    ram_cell[     497] = 32'h1d21b314;
    ram_cell[     498] = 32'h24e47509;
    ram_cell[     499] = 32'hce85ce90;
    ram_cell[     500] = 32'h4c312dbd;
    ram_cell[     501] = 32'h46b8a911;
    ram_cell[     502] = 32'h69f62744;
    ram_cell[     503] = 32'h2b28c50d;
    ram_cell[     504] = 32'h141e0826;
    ram_cell[     505] = 32'h94e739d5;
    ram_cell[     506] = 32'h990d1b18;
    ram_cell[     507] = 32'hf888d17b;
    ram_cell[     508] = 32'h8a110365;
    ram_cell[     509] = 32'ha4dbd4cc;
    ram_cell[     510] = 32'h1179aed6;
    ram_cell[     511] = 32'h18be10d9;
    // src matrix B
    ram_cell[     512] = 32'h00015f47;
    ram_cell[     513] = 32'h54092dec;
    ram_cell[     514] = 32'h0cf36a4e;
    ram_cell[     515] = 32'hb40055ba;
    ram_cell[     516] = 32'h544f9d12;
    ram_cell[     517] = 32'h8c0d806f;
    ram_cell[     518] = 32'h34ba44d2;
    ram_cell[     519] = 32'h75717e75;
    ram_cell[     520] = 32'h3ef86909;
    ram_cell[     521] = 32'hd5a9bc8b;
    ram_cell[     522] = 32'hec88f0a6;
    ram_cell[     523] = 32'h78a7e77b;
    ram_cell[     524] = 32'h7aca8a1e;
    ram_cell[     525] = 32'hd6b0f872;
    ram_cell[     526] = 32'hf5096db0;
    ram_cell[     527] = 32'hdc9c982d;
    ram_cell[     528] = 32'h71d81bbe;
    ram_cell[     529] = 32'he57a0a48;
    ram_cell[     530] = 32'h4aa42f23;
    ram_cell[     531] = 32'hb45db747;
    ram_cell[     532] = 32'h02658f51;
    ram_cell[     533] = 32'h9ae17a97;
    ram_cell[     534] = 32'h4ad4cc15;
    ram_cell[     535] = 32'hb9d98e9c;
    ram_cell[     536] = 32'h025805b6;
    ram_cell[     537] = 32'hf95039aa;
    ram_cell[     538] = 32'he37c4ead;
    ram_cell[     539] = 32'h39319641;
    ram_cell[     540] = 32'h5146f998;
    ram_cell[     541] = 32'h46408f24;
    ram_cell[     542] = 32'h239bacd4;
    ram_cell[     543] = 32'hef02eb1d;
    ram_cell[     544] = 32'hea8dec7d;
    ram_cell[     545] = 32'h8410aedf;
    ram_cell[     546] = 32'h00d830e2;
    ram_cell[     547] = 32'h48635076;
    ram_cell[     548] = 32'he9def2af;
    ram_cell[     549] = 32'hde67c152;
    ram_cell[     550] = 32'h08c81b48;
    ram_cell[     551] = 32'h4706d9b9;
    ram_cell[     552] = 32'h98d6434a;
    ram_cell[     553] = 32'h4d8ffcfe;
    ram_cell[     554] = 32'h75d3629d;
    ram_cell[     555] = 32'hde3a52a6;
    ram_cell[     556] = 32'h3549837d;
    ram_cell[     557] = 32'h4bd1523a;
    ram_cell[     558] = 32'hd3a7fab3;
    ram_cell[     559] = 32'h7ae98de4;
    ram_cell[     560] = 32'haa4e7abe;
    ram_cell[     561] = 32'hd8fd1a37;
    ram_cell[     562] = 32'hf4d1791b;
    ram_cell[     563] = 32'h3af3ec5f;
    ram_cell[     564] = 32'hcbbb0588;
    ram_cell[     565] = 32'h0f3fe247;
    ram_cell[     566] = 32'h900c568f;
    ram_cell[     567] = 32'hd8d7812a;
    ram_cell[     568] = 32'ha5f559fb;
    ram_cell[     569] = 32'hbe97ce6f;
    ram_cell[     570] = 32'h35e6534c;
    ram_cell[     571] = 32'h8179aa12;
    ram_cell[     572] = 32'h17876469;
    ram_cell[     573] = 32'he7f20401;
    ram_cell[     574] = 32'h54c7bcbf;
    ram_cell[     575] = 32'hc701d439;
    ram_cell[     576] = 32'he9e0ed6a;
    ram_cell[     577] = 32'ha78ef122;
    ram_cell[     578] = 32'hf0e90604;
    ram_cell[     579] = 32'hbda6a8df;
    ram_cell[     580] = 32'h9c5a3216;
    ram_cell[     581] = 32'hb031cba4;
    ram_cell[     582] = 32'hb39cf2c2;
    ram_cell[     583] = 32'ha859b816;
    ram_cell[     584] = 32'h5c38a817;
    ram_cell[     585] = 32'ha2a14d65;
    ram_cell[     586] = 32'h66c91371;
    ram_cell[     587] = 32'hfbc4c341;
    ram_cell[     588] = 32'h9fe35720;
    ram_cell[     589] = 32'hb497eeb2;
    ram_cell[     590] = 32'ha46b6277;
    ram_cell[     591] = 32'h38fa8985;
    ram_cell[     592] = 32'ha04dfde9;
    ram_cell[     593] = 32'h1199c8b7;
    ram_cell[     594] = 32'h28ee7f9c;
    ram_cell[     595] = 32'h1243b7ab;
    ram_cell[     596] = 32'h83f7723d;
    ram_cell[     597] = 32'h77b9eb96;
    ram_cell[     598] = 32'h0295862a;
    ram_cell[     599] = 32'h745071b6;
    ram_cell[     600] = 32'hc49d22c3;
    ram_cell[     601] = 32'h01387874;
    ram_cell[     602] = 32'h96dd5d6b;
    ram_cell[     603] = 32'h3b7cb47d;
    ram_cell[     604] = 32'hee58e390;
    ram_cell[     605] = 32'h0393ccf2;
    ram_cell[     606] = 32'hef3a6204;
    ram_cell[     607] = 32'h735bec58;
    ram_cell[     608] = 32'h34a61a76;
    ram_cell[     609] = 32'hacf7f249;
    ram_cell[     610] = 32'hfce2d5c5;
    ram_cell[     611] = 32'hcf46de12;
    ram_cell[     612] = 32'h5ff0b47b;
    ram_cell[     613] = 32'hce44a9ea;
    ram_cell[     614] = 32'h4a5cd743;
    ram_cell[     615] = 32'ha3403aed;
    ram_cell[     616] = 32'h35709c9c;
    ram_cell[     617] = 32'h650ea984;
    ram_cell[     618] = 32'ha97429f4;
    ram_cell[     619] = 32'h601797bb;
    ram_cell[     620] = 32'hd133d7d6;
    ram_cell[     621] = 32'h9be7aaef;
    ram_cell[     622] = 32'h983759da;
    ram_cell[     623] = 32'h781df2fd;
    ram_cell[     624] = 32'h9dc64c78;
    ram_cell[     625] = 32'h870cca4f;
    ram_cell[     626] = 32'ha0206205;
    ram_cell[     627] = 32'h29b558bd;
    ram_cell[     628] = 32'h1da18409;
    ram_cell[     629] = 32'h85dccef0;
    ram_cell[     630] = 32'h806ae0da;
    ram_cell[     631] = 32'h5924f5b1;
    ram_cell[     632] = 32'hf8ef95d9;
    ram_cell[     633] = 32'h96bef0df;
    ram_cell[     634] = 32'h09425ae9;
    ram_cell[     635] = 32'hb1fefc19;
    ram_cell[     636] = 32'h4ac6749f;
    ram_cell[     637] = 32'hfd5b1e92;
    ram_cell[     638] = 32'h18ad1352;
    ram_cell[     639] = 32'h97d66b20;
    ram_cell[     640] = 32'h71f6e6c5;
    ram_cell[     641] = 32'hd63bcb5e;
    ram_cell[     642] = 32'h2990b70f;
    ram_cell[     643] = 32'h30f3faf0;
    ram_cell[     644] = 32'ha4f187a2;
    ram_cell[     645] = 32'ha2d69401;
    ram_cell[     646] = 32'hb6b15550;
    ram_cell[     647] = 32'hb32061aa;
    ram_cell[     648] = 32'h58333279;
    ram_cell[     649] = 32'he8eb3f64;
    ram_cell[     650] = 32'h4c6170ff;
    ram_cell[     651] = 32'h869cc3f9;
    ram_cell[     652] = 32'hf9f29afb;
    ram_cell[     653] = 32'h4ffe7c27;
    ram_cell[     654] = 32'h4f411eef;
    ram_cell[     655] = 32'h132f93d0;
    ram_cell[     656] = 32'haae11e04;
    ram_cell[     657] = 32'h3ef6168a;
    ram_cell[     658] = 32'hd9872ca6;
    ram_cell[     659] = 32'hf720bdfd;
    ram_cell[     660] = 32'h7047a507;
    ram_cell[     661] = 32'h6e8a41f2;
    ram_cell[     662] = 32'h5bd6b773;
    ram_cell[     663] = 32'h3b3306f6;
    ram_cell[     664] = 32'h74bd4c59;
    ram_cell[     665] = 32'h6b12ebd7;
    ram_cell[     666] = 32'h52aa2f46;
    ram_cell[     667] = 32'hee38a288;
    ram_cell[     668] = 32'h2d44a978;
    ram_cell[     669] = 32'haa8ef9da;
    ram_cell[     670] = 32'h0f36cabd;
    ram_cell[     671] = 32'h19e91142;
    ram_cell[     672] = 32'h7d8455c7;
    ram_cell[     673] = 32'h07eb7f19;
    ram_cell[     674] = 32'hf777c341;
    ram_cell[     675] = 32'hcbd4257c;
    ram_cell[     676] = 32'h15becaf0;
    ram_cell[     677] = 32'hecada651;
    ram_cell[     678] = 32'h73461d54;
    ram_cell[     679] = 32'h516440ff;
    ram_cell[     680] = 32'hf73dbcd5;
    ram_cell[     681] = 32'h17ea2f05;
    ram_cell[     682] = 32'h48ab3615;
    ram_cell[     683] = 32'hd3749247;
    ram_cell[     684] = 32'h8bf7115a;
    ram_cell[     685] = 32'hb1b06d47;
    ram_cell[     686] = 32'h439881de;
    ram_cell[     687] = 32'hc4e59195;
    ram_cell[     688] = 32'h9306fb70;
    ram_cell[     689] = 32'h412f732d;
    ram_cell[     690] = 32'hc1744386;
    ram_cell[     691] = 32'h03f958e1;
    ram_cell[     692] = 32'he51b84ff;
    ram_cell[     693] = 32'hc6ec14ee;
    ram_cell[     694] = 32'h65ec85d2;
    ram_cell[     695] = 32'he49f0672;
    ram_cell[     696] = 32'h787205bc;
    ram_cell[     697] = 32'hfd02cecc;
    ram_cell[     698] = 32'h13e9afb2;
    ram_cell[     699] = 32'hd5061d02;
    ram_cell[     700] = 32'hb635d535;
    ram_cell[     701] = 32'hd8c292e9;
    ram_cell[     702] = 32'hdb405533;
    ram_cell[     703] = 32'hfe920a0e;
    ram_cell[     704] = 32'h7937def6;
    ram_cell[     705] = 32'hb5d225e0;
    ram_cell[     706] = 32'hb165f9ab;
    ram_cell[     707] = 32'h3036c089;
    ram_cell[     708] = 32'hf05313a2;
    ram_cell[     709] = 32'h3d4a649d;
    ram_cell[     710] = 32'hd7e5b692;
    ram_cell[     711] = 32'h00d16ac7;
    ram_cell[     712] = 32'h2820c68b;
    ram_cell[     713] = 32'h21cfc66d;
    ram_cell[     714] = 32'h7dce968c;
    ram_cell[     715] = 32'he1dbb201;
    ram_cell[     716] = 32'h0e7e12bb;
    ram_cell[     717] = 32'h8f643654;
    ram_cell[     718] = 32'he4b38f75;
    ram_cell[     719] = 32'h477189fd;
    ram_cell[     720] = 32'hb71baeb0;
    ram_cell[     721] = 32'h3f2d50a6;
    ram_cell[     722] = 32'hfe4f2554;
    ram_cell[     723] = 32'h4f151c76;
    ram_cell[     724] = 32'h2af9503b;
    ram_cell[     725] = 32'h94aa7201;
    ram_cell[     726] = 32'heff3e6fc;
    ram_cell[     727] = 32'he513ff78;
    ram_cell[     728] = 32'h3d673010;
    ram_cell[     729] = 32'ha4d9c8a7;
    ram_cell[     730] = 32'hf13e9b8d;
    ram_cell[     731] = 32'h4bb3f0a8;
    ram_cell[     732] = 32'h712b0ef0;
    ram_cell[     733] = 32'h9faf6296;
    ram_cell[     734] = 32'h3aa2e1f1;
    ram_cell[     735] = 32'hf0d6c217;
    ram_cell[     736] = 32'h4297971e;
    ram_cell[     737] = 32'h1bc1078b;
    ram_cell[     738] = 32'hcc5b0dbe;
    ram_cell[     739] = 32'h97f21acc;
    ram_cell[     740] = 32'h3ea44de5;
    ram_cell[     741] = 32'h0b7ed373;
    ram_cell[     742] = 32'h749a4348;
    ram_cell[     743] = 32'h04994e79;
    ram_cell[     744] = 32'h6d0bfaf3;
    ram_cell[     745] = 32'h66436b31;
    ram_cell[     746] = 32'h694bd69b;
    ram_cell[     747] = 32'h17f48d13;
    ram_cell[     748] = 32'hc93edd62;
    ram_cell[     749] = 32'h25f8fa5f;
    ram_cell[     750] = 32'hd3cd30d0;
    ram_cell[     751] = 32'hf9e91671;
    ram_cell[     752] = 32'h5b9a281c;
    ram_cell[     753] = 32'hf206a596;
    ram_cell[     754] = 32'h89caad13;
    ram_cell[     755] = 32'hf126755d;
    ram_cell[     756] = 32'h500199ed;
    ram_cell[     757] = 32'hdb6883d1;
    ram_cell[     758] = 32'h0a26b40b;
    ram_cell[     759] = 32'h470f1672;
    ram_cell[     760] = 32'h7e064dc5;
    ram_cell[     761] = 32'hbc0b4fcc;
    ram_cell[     762] = 32'hc34e59f3;
    ram_cell[     763] = 32'h352d538b;
    ram_cell[     764] = 32'hc88f6111;
    ram_cell[     765] = 32'h2b0ba254;
    ram_cell[     766] = 32'h646be84a;
    ram_cell[     767] = 32'h6cbab852;
end

endmodule

